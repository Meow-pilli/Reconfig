// sincos.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
/*
module sincos (
		input  wire [9:0] a,      //      a.a
		input  wire       areset, // areset.reset
		output wire [4:0] c,      //      c.c
		input  wire       clk,    //    clk.clk
		output wire [4:0] s       //      s.s
	);

	sincos_CORDIC_0 cordic_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.a      (a),      //      a.a
		.c      (c),      //      c.c
		.s      (s)       //      s.s
	);

endmodule
*/

module sincos(
	input [9:0]a,
	input areset,
	input clk,
	output [6:0]sin_sev_dec, // sin decimal
	output [6:0]sin_sev_int, // sin integer
	output [6:0]sin_sev_sign, // sin sign
	output [6:0]cos_sev_dec, // cos decimal
	output [6:0]cos_sev_int, // cos integer
	output [6:0]cos_sev_sign  // ocs sign
	);

	reg [4:0]temp_cos;
	reg [4:0]temp_sin;

	sincos_CORDIC_0 u0(.a(a), .areset(!areset), .clk(clk), .c(temp1), .s(temp2)); 
	seven_display_decoder u1(.in(temp_cos[2:0]), .out(cos_sev_dec));
	seven_display_decoder u2(.in(temp_cos[3]), .out(cos_sev_int));
	seven_display_decoder u3(.in(temp_cos[4]), .out(cos_sev_sign));
	seven_display_decoder u4(.in(temp_sin[2:0]), .out(sin_sev_dec));
	seven_display_decoder u5(.in(temp_sin[3]), .out(sin_sev_int));
	seven_display_decoder u6(.in(temp_sin[4]), .out(sin_sev_sign));

endmodule

module seven_display_decoder(
	input wire [2:0]in,
	output reg [6:0]out
);
always @(*) begin
    case(in)
        3'b000: out = 7'b1000000; // Display 0
        3'b001: out = 7'b1111001; // Display 1
        3'b010: out = 7'b0100100; // Display 2
        3'b011: out = 7'b0110000; // Display 3
        3'b100: out = 7'b0011001; // Display 4
        3'b101: out = 7'b0010010; // Display 5
        3'b110: out = 7'b0000010; // Display 6
        3'b111: out = 7'b1111000; // Display 7
        default: out = 7'b1111111; // Turn off all segments for unknown input
    endcase
end
endmodule
/*
module seven_display_decoder(
	input wire in,
	output reg [6:0]out
);
always @(*) begin
    case(in)
        3'b000: out = 7'b1000000; // Display 0
        3'b001: out = 7'b1111001; // Display 1
        3'b010: out = 7'b0100100; // Display 2
        3'b011: out = 7'b0110000; // Display 3
        3'b100: out = 7'b0011001; // Display 4
        3'b101: out = 7'b0010010; // Display 5
        3'b110: out = 7'b0000010; // Display 6
        3'b111: out = 7'b1111000; // Display 7
        default: out = 7'b1111111; // Turn off all segments for unknown input
    endcase
end
endmodule
*/