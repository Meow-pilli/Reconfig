
module sincos (
	clk,
	areset,
	a,
	c,
	s);	

	input		clk;
	input		areset;
	input	[9:0]	a;
	output	[2:0]	c;
	output	[2:0]	s;
endmodule
